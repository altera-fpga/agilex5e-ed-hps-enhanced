// Copyright (C) 2021 Intel Corporation.
// SPDX-License-Identifier: MIT

//
// Description
//-----------------------------------------------------------------------------
//
// This package defines the global parameters of FIM
//
//----------------------------------------------------------------------------

`ifndef __OFS_FIM_CFG_PKG_SV__
`define __OFS_FIM_CFG_PKG_SV__

// IP configuration database, generated by OFS script ofs_ip_cfg_db.tcl after
// IP generation.
//`include "ofs_ip_cfg_db.vh"
//
// Generated by OFS script iopll_get_cfg.tcl using qsys-script
//

`ifndef __OFS_FIM_IP_CFG_SYS_CLK__
`define __OFS_FIM_IP_CFG_SYS_CLK__ 1

//
// Clock frequencies and names
//
`define OFS_FIM_IP_CFG_SYS_CLK_CLK0_NAME     clk_sys
`define OFS_FIM_IP_CFG_SYS_CLK_CLK0_MHZ      470.0
`define OFS_FIM_IP_CFG_SYS_CLK_CLK0_MHZ_INT  470  // Nearest integer frequency

`define OFS_FIM_IP_CFG_SYS_CLK_CLK1_NAME     clk_100m
`define OFS_FIM_IP_CFG_SYS_CLK_CLK1_MHZ      100.0
`define OFS_FIM_IP_CFG_SYS_CLK_CLK1_MHZ_INT  100  // Nearest integer frequency

`define OFS_FIM_IP_CFG_SYS_CLK_CLK2_NAME     clk_sys_div2
`define OFS_FIM_IP_CFG_SYS_CLK_CLK2_MHZ      235.0
`define OFS_FIM_IP_CFG_SYS_CLK_CLK2_MHZ_INT  235  // Nearest integer frequency

`define OFS_FIM_IP_CFG_SYS_CLK_CLK3_NAME     clk_ptp_slv
`define OFS_FIM_IP_CFG_SYS_CLK_CLK3_MHZ      155.555556
`define OFS_FIM_IP_CFG_SYS_CLK_CLK3_MHZ_INT  156  // Nearest integer frequency

`define OFS_FIM_IP_CFG_SYS_CLK_CLK4_NAME     clk_50m
`define OFS_FIM_IP_CFG_SYS_CLK_CLK4_MHZ      50.0
`define OFS_FIM_IP_CFG_SYS_CLK_CLK4_MHZ_INT  50  // Nearest integer frequency

`define OFS_FIM_IP_CFG_SYS_CLK_CLK5_NAME     clk_sys_div4
`define OFS_FIM_IP_CFG_SYS_CLK_CLK5_MHZ      117.5
`define OFS_FIM_IP_CFG_SYS_CLK_CLK5_MHZ_INT  118  // Nearest integer frequency

`endif // `ifndef __OFS_FIM_IP_CFG_SYS_CLK__
//
// Generated by OFS script pcie_ss_get_cfg.tcl using qsys-script
//

`ifndef __OFS_FIM_IP_CFG_PCIE_SS__
`define __OFS_FIM_IP_CFG_PCIE_SS__ 1

//
// The OFS_FIM_IP_CFG_<ip_name>_PF<n>_ACTIVE macro will be defined iff the
// PF is active. The value does not have to be tested.
//
// For each active PF<n>, OFS_FIM_IP_CFG_<ip_name>_PF<n>_NUM_VFS will be
// defined iff there are VFs associated with the PF.
//
`define OFS_FIM_IP_CFG_PCIE_SS_PF0_ACTIVE 1
`define OFS_FIM_IP_CFG_PCIE_SS_PF0_BAR0_ADDR_WIDTH 21

`define OFS_FIM_IP_CFG_PCIE_SS_PF1_ACTIVE 1
`define OFS_FIM_IP_CFG_PCIE_SS_PF1_BAR0_ADDR_WIDTH 12


//
// The macros below represent the raw PF/VF configuration above in
// ways that are easier to process in SystemVerilog loops.
//

// Total number of PFs, not necessarily dense (see MAX_PF_NUM)
`define OFS_FIM_IP_CFG_PCIE_SS_NUM_PFS 2
// Total number of VFs across all PFs
`define OFS_FIM_IP_CFG_PCIE_SS_TOTAL_NUM_VFS 0
// Largest active PF number
`define OFS_FIM_IP_CFG_PCIE_SS_MAX_PF_NUM 1
// Largest number of VFs associated with a single PF
`define OFS_FIM_IP_CFG_PCIE_SS_MAX_VFS_PER_PF 0

// Vector indicating enabled PFs (1 if enabled) with
// index range 0 to OFS_FIM_IP_CFG_PCIE_SS_MAX_PF_NUM
`define OFS_FIM_IP_CFG_PCIE_SS_PF_ENABLED_VEC 1, 1
// Vector with the number of VFs indexed by PF
`define OFS_FIM_IP_CFG_PCIE_SS_NUM_VFS_VEC 0, 0


`endif // `ifndef __OFS_FIM_IP_CFG_PCIE_SS__
//
// Generated by OFS script pcie_ss_get_cfg.tcl using qsys-script
//

`ifndef __OFS_FIM_IP_CFG_SOC_PCIE_SS__
`define __OFS_FIM_IP_CFG_SOC_PCIE_SS__ 1

//
// The OFS_FIM_IP_CFG_<ip_name>_PF<n>_ACTIVE macro will be defined iff the
// PF is active. The value does not have to be tested.
//
// For each active PF<n>, OFS_FIM_IP_CFG_<ip_name>_PF<n>_NUM_VFS will be
// defined iff there are VFs associated with the PF.
//
`define OFS_FIM_IP_CFG_SOC_PCIE_SS_PF0_ACTIVE 1
`define OFS_FIM_IP_CFG_SOC_PCIE_SS_PF0_BAR0_ADDR_WIDTH 21
`define OFS_FIM_IP_CFG_SOC_PCIE_SS_PF0_NUM_VFS 3
`define OFS_FIM_IP_CFG_SOC_PCIE_SS_PF0_VF_BAR0_ADDR_WIDTH 21


//
// The macros below represent the raw PF/VF configuration above in
// ways that are easier to process in SystemVerilog loops.
//

// Total number of PFs, not necessarily dense (see MAX_PF_NUM)
`define OFS_FIM_IP_CFG_SOC_PCIE_SS_NUM_PFS 1
// Total number of VFs across all PFs
`define OFS_FIM_IP_CFG_SOC_PCIE_SS_TOTAL_NUM_VFS 3
// Largest active PF number
`define OFS_FIM_IP_CFG_SOC_PCIE_SS_MAX_PF_NUM 0
// Largest number of VFs associated with a single PF
`define OFS_FIM_IP_CFG_SOC_PCIE_SS_MAX_VFS_PER_PF 3

// Vector indicating enabled PFs (1 if enabled) with
// index range 0 to OFS_FIM_IP_CFG_SOC_PCIE_SS_MAX_PF_NUM
`define OFS_FIM_IP_CFG_SOC_PCIE_SS_PF_ENABLED_VEC 1
// Vector with the number of VFs indexed by PF
`define OFS_FIM_IP_CFG_SOC_PCIE_SS_NUM_VFS_VEC 3


`endif // `ifndef __OFS_FIM_IP_CFG_SOC_PCIE_SS__
//
// Generated by OFS script hssi_ss_get_cfg.tcl using qsys-script
//

`ifndef __OFS_FIM_IP_CFG_HSSI_SS__
`define __OFS_FIM_IP_CFG_HSSI_SS__ 1

//
// The OFS_FIM_IP_CFG_<ip_name>_ETH_PORTS macro will be defined iff the
// port is active. The value does not have to be tested.
//

//
// The macros below represent the raw eth port configuration above in
// ways that are easier to process in SystemVerilog loops.
//

`define ETH_100G


`define INST_ALL_PORTS \
   `HSSI_PORT_INST(0) \
   `HSSI_PORT_INST(4) \


`define INCLUDE_HSSI_PORT_0
`define INCLUDE_HSSI_PORT_4

`define ENUM_PORT_INDEX PORT_0, PORT_4,


`define INST_ALL_LED_0(led_type, led_idx, operator) \
    `INST_LED(``led_type``,0,``led_idx``, operator) \

`define INST_ALL_LED_1(led_type, led_idx, operator) \
    `INST_LED(``led_type``,4,``led_idx``, operator) \


// Total number of ports, not necessarily dense (see MAX_PORT_NUM)
`define OFS_FIM_IP_CFG_HSSI_SS_NUM_ETH_PORTS 2
`define OFS_FIM_IP_CFG_HSSI_SS_ETH_PACKET_WIDTH 512
`define OFS_FIM_IP_CFG_HSSI_SS_NUM_LANES 4


`endif // `ifndef __OFS_FIM_IP_CFG_HSSI_SS__
//
// Generated by OFS script mem_ss_get_cfg.tcl using qsys-script
//

`ifndef __OFS_FIM_IP_CFG_MEM_SS__
`define __OFS_FIM_IP_CFG_MEM_SS__ 1


//
// Flags to enable memory channel instantiation/configuration
//
`define OFS_FIM_IP_CFG_MEM_SS_EN_MEM_3
`define OFS_FIM_IP_CFG_MEM_SS_EN_MEM_2
`define OFS_FIM_IP_CFG_MEM_SS_EN_MEM_1
`define OFS_FIM_IP_CFG_MEM_SS_EN_MEM_0
`define OFS_FIM_IP_CFG_MEM_SS_NUM_MEM_CHANNELS 4

//
// AXI-MM user interface configuration
//
`define OFS_FIM_IP_CFG_MEM_SS_DEFINES_USER_AXI 1
`define OFS_FIM_IP_CFG_MEM_SS_AXI_DATA_WIDTH 512
`define OFS_FIM_IP_CFG_MEM_SS_AXI_USER_WIDTH 1
`define OFS_FIM_IP_CFG_MEM_SS_AXI_LEN_WIDTH 8
`define OFS_FIM_IP_CFG_MEM_SS_AXI_ID_WIDTH 9
`define OFS_FIM_IP_CFG_MEM_SS_AXI_ADDR_WIDTH 32

//
// Fabric EMIF interface configuration
//
`define OFS_FIM_IP_CFG_MEM_SS_DEFINES_EMIF_DDR4 1
`define OFS_FIM_IP_CFG_MEM_SS_DDR4_A_WIDTH 17
`define OFS_FIM_IP_CFG_MEM_SS_DDR4_BA_WIDTH 2
`define OFS_FIM_IP_CFG_MEM_SS_DDR4_BG_WIDTH 1
`define OFS_FIM_IP_CFG_MEM_SS_DDR4_CK_WIDTH 1
`define OFS_FIM_IP_CFG_MEM_SS_DDR4_CKE_WIDTH 1
`define OFS_FIM_IP_CFG_MEM_SS_DDR4_CS_N_WIDTH 1
`define OFS_FIM_IP_CFG_MEM_SS_DDR4_ODT_WIDTH 1
`define OFS_FIM_IP_CFG_MEM_SS_DDR4_DQ_WIDTH 32

`endif // `ifndef __OFS_FIM_IP_CFG_MEM_SS__
package ofs_fim_cfg_pkg;

localparam MAIN_CLK_MHZ = `OFS_FIM_IP_CFG_SYS_CLK_CLK0_MHZ_INT;

//*****************
// PCIe host parameters
//*****************
`ifdef SIM_USE_PCIE_GEN3X16_BFM
   localparam PCIE_LANES = 16;
`else
   localparam PCIE_LANES = 16;
`endif

localparam NUM_PCIE_HOST      = 1;
localparam PCIE_HOST_WIDTH    = $clog2(NUM_PCIE_HOST);

localparam PCIE_TDATA_WIDTH  = 512;
localparam PCIE_TUSER_WIDTH  = 10;
localparam PCIE_LITE_CSR_WIDTH = 20;

localparam PCIE_RP_MAX_TAGS   = (1<<10);
localparam PCIE_RP_TAG_WIDTH  = $clog2(PCIE_RP_MAX_TAGS);

localparam MAX_PAYLOAD_SIZE   = 128; // DW
localparam MAX_RD_REQ_SIZE    = 128; // DW

//*****************
// MMIO parameters
//*****************
localparam PORTS              = 1;
localparam MMIO_TID_WIDTH     = PCIE_HOST_WIDTH + PCIE_RP_TAG_WIDTH; // Matches PCIe TLP tag width
localparam MMIO_DATA_WIDTH    = 64;
localparam MMIO_ADDR_WIDTH    = `OFS_FIM_IP_CFG_SOC_PCIE_SS_PF0_BAR0_ADDR_WIDTH;

//MSIX
`ifdef NUM_AFUS
localparam   NUM_AFUS    = 2;
`else
localparam   NUM_AFUS    = 1;
`endif
localparam LNUM_AFUS = NUM_AFUS>1?$clog2(NUM_AFUS):1'h1;
localparam NUM_AFU_INTERRUPTS = 7;
localparam L_NUM_AFU_INTERRUPTS = $clog2(NUM_AFU_INTERRUPTS);


endpackage

`endif // __OFS_FIM_CFG_PKG_SV__
