module pv_ss_mem_msa_tg
  #(
    parameter ADDR_WIDTH      = 31,
    parameter DATA_WIDTH      = 256,
    parameter ID_W_WIDTH      = 9,
    parameter ID_R_WIDTH      = 9,
    parameter USER_REQ_WIDTH  = 1,
    parameter USER_RESP_WIDTH = 1,
    parameter USER_DATA_WIDTH = 1
    )
  (
   input wire                        ninit_done,
   output wire                       traffic_gen_pass,
   output wire                       traffic_gen_fail,
   output wire                       traffic_gen_timeout,
   input wire [19:0]                 tg_cfg_address,
   input wire                        tg_cfg_write,
   input wire [31:0]                 tg_cfg_writedata,
   input wire                        tg_cfg_read,
   output wire [31:0]                tg_cfg_readdata,
   output wire                       tg_cfg_readdatavalid,
   output wire                       tg_cfg_waitrequest,
   output wire [ID_W_WIDTH-1:0]      axi_awid,
   output wire [ADDR_WIDTH-1:0]      axi_awaddr,
   output wire                       axi_awvalid,
   output wire [0:0]                 axi_awuser,
   output wire [7:0]                 axi_awlen,
   output wire [2:0]                 axi_awsize,
   output wire [1:0]                 axi_awburst,
   input wire                        axi_awready,
   output wire [0:0]                 axi_awlock,
   output wire [3:0]                 axi_awcache,
   output wire [2:0]                 axi_awprot,
   output wire [ID_R_WIDTH-1:0]      axi_arid,
   output wire [ADDR_WIDTH-1:0]      axi_araddr,
   output wire                       axi_arvalid,
   output wire [USER_REQ_WIDTH-1:0]  axi_aruser,
   output wire [7:0]                 axi_arlen,
   output wire [2:0]                 axi_arsize,
   output wire [1:0]                 axi_arburst,
   input wire                        axi_arready,
   output wire [0:0]                 axi_arlock,
   output wire [3:0]                 axi_arcache,
   output wire [2:0]                 axi_arprot,
   output wire [DATA_WIDTH-1:0]      axi_wdata,
   output wire [USER_DATA_WIDTH-1:0] axi_wuser,
   output wire [DATA_WIDTH/8-1:0]    axi_wstrb,
   output wire                       axi_wlast,
   output wire                       axi_wvalid,
   input wire                        axi_wready,
   input wire [ID_W_WIDTH-1:0]       axi_bid,
   input wire [1:0]                  axi_bresp,
   input wire [USER_RESP_WIDTH-1:0]  axi_buser,
   input wire                        axi_bvalid,
   output wire                       axi_bready,
   input wire [DATA_WIDTH-1:0]       axi_rdata,
   input wire [1:0]                  axi_rresp,
   input wire [USER_RESP_WIDTH-1:0]  axi_ruser,
   input wire                        axi_rlast,
   input wire                        axi_rvalid,
   output wire                       axi_rready,
   input wire [ID_R_WIDTH-1:0]       axi_rid,
   input wire                        emif_usr_clk,
   input wire                        emif_usr_reset_n
   );

   localparam WORD_ADDR_WIDTH = ADDR_WIDTH - $clog2(DATA_WIDTH/8);


   altera_emif_avl_tg_2_top
     #(
       .PROTOCOL_ENUM                         ("PROTOCOL_DDR4"),
       .BYPASS_DEFAULT_PATTERN                (1),
       .BYPASS_USER_STAGE                     (0),
       .USE_AVL_BYTEEN                        (0),
       .AMM_WORD_ADDRESS_WIDTH                (WORD_ADDR_WIDTH),
       .PORT_TG_CFG_ADDRESS_WIDTH             (10),
       .PORT_TG_CFG_RDATA_WIDTH               (32),
       .PORT_TG_CFG_WDATA_WIDTH               (32),
       .DIAG_EXPORT_TG_CFG_AVALON_SLAVE       ("TG_CFG_AMM_EXPORT_MODE_EXPORT"),
       .MEM_TTL_DATA_WIDTH                    (32),
       .MEM_TTL_NUM_OF_WRITE_GROUPS           (4),
       .AVL_TO_DQ_WIDTH_RATIO                 (8),
       .CTRL_INTERFACE_TYPE                   ("AXI"),
       .PORT_CTRL_AXI4_AWID_WIDTH             (ID_W_WIDTH),
       .PORT_CTRL_AXI4_AWADDR_WIDTH           (ADDR_WIDTH),
       .PORT_CTRL_AXI4_AWUSER_WIDTH           (USER_REQ_WIDTH),
       .PORT_CTRL_AXI4_AWLEN_WIDTH            (8),
       .PORT_CTRL_AXI4_AWSIZE_WIDTH           (3),
       .PORT_CTRL_AXI4_AWBURST_WIDTH          (2),
       .PORT_CTRL_AXI4_AWLOCK_WIDTH           (1),
       .PORT_CTRL_AXI4_AWCACHE_WIDTH          (4),
       .PORT_CTRL_AXI4_AWPROT_WIDTH           (3),
       .PORT_CTRL_AXI4_ARID_WIDTH             (ID_R_WIDTH),
       .PORT_CTRL_AXI4_ARADDR_WIDTH           (ADDR_WIDTH),
       .PORT_CTRL_AXI4_ARUSER_WIDTH           (USER_REQ_WIDTH),
       .PORT_CTRL_AXI4_ARLEN_WIDTH            (8),
       .PORT_CTRL_AXI4_ARSIZE_WIDTH           (3),
       .PORT_CTRL_AXI4_ARBURST_WIDTH          (2),
       .PORT_CTRL_AXI4_ARLOCK_WIDTH           (1),
       .PORT_CTRL_AXI4_ARCACHE_WIDTH          (4),
       .PORT_CTRL_AXI4_ARPROT_WIDTH           (3),
       .PORT_CTRL_AXI4_WDATA_WIDTH            (DATA_WIDTH),
       .PORT_CTRL_AXI4_WUSER_WIDTH            (USER_DATA_WIDTH),
       .PORT_CTRL_AXI4_WSTRB_WIDTH            (DATA_WIDTH/8),
       .PORT_CTRL_AXI4_BID_WIDTH              (ID_W_WIDTH),
       .PORT_CTRL_AXI4_BRESP_WIDTH            (2),
       .PORT_CTRL_AXI4_BUSER_WIDTH            (USER_RESP_WIDTH),
       .PORT_CTRL_AXI4_RID_WIDTH              (ID_R_WIDTH),
       .PORT_CTRL_AXI4_RDATA_WIDTH            (DATA_WIDTH),
       .PORT_CTRL_AXI4_RRESP_WIDTH            (2),
       .PORT_CTRL_AXI4_RUSER_WIDTH            (USER_RESP_WIDTH),
       .RW_RPT_COUNT_WIDTH                    (32),
       .RW_OPERATION_COUNT_WIDTH              (32),
       .RW_LOOP_COUNT_WIDTH                   (32)
       )
   tg_0
     (
      .emif_usr_reset_n                (emif_usr_reset_n),
      .ninit_done                      (ninit_done),
      .emif_usr_clk                    (emif_usr_clk),
      .axi_awid                        (axi_awid),
      .axi_awaddr                      (axi_awaddr),
      .axi_awvalid                     (axi_awvalid),
      .axi_awuser                      (axi_awuser),
      .axi_awlen                       (axi_awlen),
      .axi_awsize                      (axi_awsize),
      .axi_awburst                     (axi_awburst),
      .axi_awready                     (axi_awready),
      .axi_awlock                      (axi_awlock),
      .axi_awcache                     (axi_awcache),
      .axi_awprot                      (axi_awprot),
      .axi_arid                        (axi_arid),
      .axi_araddr                      (axi_araddr),
      .axi_arvalid                     (axi_arvalid),
      .axi_aruser                      (axi_aruser),
      .axi_arlen                       (axi_arlen),
      .axi_arsize                      (axi_arsize),
      .axi_arburst                     (axi_arburst),
      .axi_arready                     (axi_arready),
      .axi_arlock                      (axi_arlock),
      .axi_arcache                     (axi_arcache),
      .axi_arprot                      (axi_arprot),
      .axi_wdata                       (axi_wdata),
//      .axi_wuser                       (axi_wuser),
      .axi_wstrb                       (axi_wstrb),
      .axi_wlast                       (axi_wlast),
      .axi_wvalid                      (axi_wvalid),
      .axi_wready                      (axi_wready),
      .axi_bid                         (axi_bid),
      .axi_bresp                       (axi_bresp),
      .axi_buser                       (axi_buser),
      .axi_bvalid                      (axi_bvalid),
      .axi_bready                      (axi_bready),
      .axi_rdata                       (axi_rdata),
      .axi_rresp                       (axi_rresp),
      .axi_ruser                       (axi_ruser),
      .axi_rlast                       (axi_rlast),
      .axi_rvalid                      (axi_rvalid),
      .axi_rready                      (axi_rready),
      .axi_rid                         (axi_rid),
      .traffic_gen_pass                (traffic_gen_pass),
      .traffic_gen_fail                (traffic_gen_fail),
      .traffic_gen_timeout             (traffic_gen_timeout),
      .ss_base_csr_axi4l_awaddr        (),
      .ss_base_csr_axi4l_awvalid       (),
      .ss_base_csr_axi4l_awready       (1'b0),
      .ss_base_csr_axi4l_awprot        (),
      .ss_base_csr_axi4l_araddr        (),
      .ss_base_csr_axi4l_arvalid       (),
      .ss_base_csr_axi4l_arready       (1'b0),
      .ss_base_csr_axi4l_arprot        (),
      .ss_base_csr_axi4l_wdata         (),
      .ss_base_csr_axi4l_wstrb         (),
      .ss_base_csr_axi4l_wvalid        (),
      .ss_base_csr_axi4l_wready        (1'b0),
      .ss_base_csr_axi4l_bresp         (2'b00),
      .ss_base_csr_axi4l_bvalid        (1'b0),
      .ss_base_csr_axi4l_bready        (),
      .ss_base_csr_axi4l_rdata         (32'b00000000000000000000000000000000),
      .ss_base_csr_axi4l_rresp         (2'b00),
      .ss_base_csr_axi4l_rvalid        (1'b0),
      .ss_base_csr_axi4l_rready        (),
      .ctrl_user_priority_hi_0         (),
      .ctrl_auto_precharge_req_0       (),
      .ctrl_ecc_user_interrupt_0       (1'b0),
      .ctrl_ecc_readdataerror_0        (1'b0),
      .mmr_master_waitrequest_0        (1'b0),
      .mmr_master_read_0               (),
      .mmr_master_write_0              (),
      .mmr_master_address_0            (),
      .mmr_master_readdata_0           (32'b00000000000000000000000000000000),
      .mmr_master_writedata_0          (),
      .mmr_master_burstcount_0         (),
      .mmr_master_beginbursttransfer_0 (),
      .mmr_master_readdatavalid_0      (1'b0),

      // ***** START CHANGE *****
      .tg_cfg_waitrequest              (tg_cfg_waitrequest),
      .tg_cfg_read                     (tg_cfg_read),
      .tg_cfg_write                    (tg_cfg_write),
      .tg_cfg_address                  (tg_cfg_address[9:0]),
      .tg_cfg_readdata                 (tg_cfg_readdata),
      .tg_cfg_writedata                (tg_cfg_writedata),
      .tg_cfg_readdatavalid            (tg_cfg_readdatavalid)
      // ***** END CHANGE *****
      );

endmodule
