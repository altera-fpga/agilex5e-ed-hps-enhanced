// Copyright (C) 2021 Intel Corporation.
// SPDX-License-Identifier: MIT

`ifndef fpga_defines
	`define fpga_defines

   //--------------------------------------------------------------------
   //  Technology
   //--------------------------------------------------------------------
   `define FAMILY  "Agilex" // Targeted Device Family
   `define DEVICE_FAMILY  "Agilex" // Targeted Device Family
   `define DEVICE_FAMILY_IS_AGILEX
   `define PTILE
   `define ETILE
 `endif
